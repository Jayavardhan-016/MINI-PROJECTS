module tb;
  reg [9:0]a,b,c;
  initial begin 
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b1111111111;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b0011000000;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b0000110000;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b0000001100;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b1111111111;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
    a=10'b1111111111;b=10'b1111111111;c=10'b1111111111;#5;
    a=10'b0000110000;b=10'b1100110011;c=10'b1100110000;#5;
    a=10'b0000110000;b=10'b1100110011;c=10'b1100110000;#5;
    a=10'b0000110000;b=10'b1100110011;c=10'b1100110000;#5;
    a=10'b1111111111;b=10'b1100110011;c=10'b1100110000;#5;
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
    a=10'b1111111111;b=10'b1111111111;c=10'b1111111111;#5;
    a=10'b1100110000;b=10'b0000000011;c=10'b1100000011;#5;
    a=10'b1100110000;b=10'b0000011111;c=10'b1100000011;#5;
    a=10'b1100110000;b=10'b0000000011;c=10'b1100000011;#5;
    a=10'b1111111111;b=10'b1111111111;c=10'b1111111111;#5;
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
    a=10'b1111111111;b=10'b1100000011;c=10'b1111111111;#5;
    a=10'b1100110000;b=10'b0011001100;c=10'b0000000011;#5;
    a=10'b1100110000;b=10'b0000110000;c=10'b0000000011;#5;
    a=10'b1100110000;b=10'b0011000000;c=10'b0000000011;#5;
    a=10'b1111110000;b=10'b1100000000;c=10'b0000000011;#5;
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
    a=10'b1111111111;b=10'b1111111111;c=10'b1111111111;#5;
    a=10'b1100110000;b=10'b1100110011;c=10'b0001111000;#5;
    a=10'b1100110000;b=10'b1100110011;c=10'b0011001100;#5;
    a=10'b1100110000;b=10'b1100110011;c=10'b0110000110;#5;
    a=10'b1111110000;b=10'b1100110011;c=10'b1100000011;#5;
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
    a=10'b1100000011;b=10'b1111111111;c=10'b1111110011;#5;
    a=10'b0011001100;b=10'b1100110000;c=10'b1100110011;#5;
    a=10'b0000110000;b=10'b1100110000;c=10'b1100110011;#5;
    a=10'b0011000000;b=10'b0110110000;c=10'b1100110011;#5;
    a=10'b1100000000;b=10'b1111111111;c=10'b1100111111;#5;
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b1111111111;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b1100111000;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b1100111100;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b1100110110;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b1111110011;c=10'b0000000000;#5;
    a=10'b0000000000;b=10'b0000000000;c=10'b0000000000;#5;
     $finish;
  end
endmodule
